library verilog;
use verilog.vl_types.all;
entity multiplicator_test is
    generic(
        data_width      : integer := 8
    );
end multiplicator_test;
